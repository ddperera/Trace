BZh91AY&SY�s� �߀Px����߰����P>rN#��k]݄�M&�OM��mM�� ����I�i��h�4h4 h4   �H)��(�4�mF�=  A�4�ɓF�� �0F`( A��F���1��  6���] � �	�`�ۼg�b&%.����&�)�`�E�t��!%`�*De��� 3(�n�6ߏQI�q�qҒ�YIҶIy��ȹP�ɖ�.�GcuZ����j�p�"$���N[�BK��+�̾"@NuJBB�=��i��Y�Ƙ��'��_�\Zv��fݳ:`���1�	��l�u�oQ���f�s׊�B%�B�Ai
�h2N�e�:4	Q
��]��a�QB
#j ��!P�2f���d$�Պ�iJg�R�,qh����5xVS�,�qe�0$sJI�3}wG;���m�$���L֠X��2�R�3Y�J�S��(�
ÉX�:]�Q*;�}l(4#����~L����.mYU������Ut$*��ɞ���xb�|�!��W0��BR�E��Oڭ�?_:&�`G�t�2��m�a���)�#yM<b��H#���� �9 "hb�������/�m���iX	�zn\���&-ش�Å&H]�zM,�+#�L��M5�du�#��\e,`~�2T!�,����l�QCl�A�K�b=����#�`Es��4j��a���b$@P���+'̺��i�"6Q��^����zP��Ɩ�ZA~��L\�:�ȵI�N`�x�a�S�4�@d��b)$��@%��	�Q�Wk���3D��/%�Qc�LH��ÓٷP����@#�H\ȳwT8��N+39Y9Èm���1�!�Q�]��$kLkv��@�Q"ɒ\�抶�M�V���@J��h��#~����	�gH��d2����g�T ��m�]t���.V�¶�L�țLO�\(n��/�촹ʝW��������(���M��rE8P��s�